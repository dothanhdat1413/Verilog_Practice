module LCD ();


endmodule